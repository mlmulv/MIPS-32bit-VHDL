library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity zero_extend is
	port (
		input : std_logic_vector(9 downto 0);
		output : std_logic_vector (31 downto 0)
	);
end zero_extend;

architecture bhv of zero_extend is 


begin

	
end bhv;